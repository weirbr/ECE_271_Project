module remote_reciever (
			input logic remote_in,
			output logic [11:0] remote_out);
			
endmodule