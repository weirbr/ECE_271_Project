module N64_reciever (
			input logic N64_in,
			output logic [11:0] N64_out);
			
endmodule